// soc_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module soc_system (
		output wire [15:0] avalon_camera_export_height,           //   avalon_camera_export.height
		output wire [15:0] avalon_camera_export_startrow,         //                       .startrow
		output wire [15:0] avalon_camera_export_startcol,         //                       .startcol
		output wire [15:0] avalon_camera_export_colmode,          //                       .colmode
		output wire [15:0] avalon_camera_export_exposure,         //                       .exposure
		output wire [15:0] avalon_camera_export_rowsize,          //                       .rowsize
		output wire [15:0] avalon_camera_export_colsize,          //                       .colsize
		output wire [15:0] avalon_camera_export_rowmode,          //                       .rowmode
		output wire        avalon_camera_export_soft_reset_n,     //                       .soft_reset_n
		output wire [15:0] avalon_camera_export_width,            //                       .width
		output wire [15:0] avalon_camera_export_h_blanking,       //                       .h_blanking
		output wire [15:0] avalon_camera_export_v_blanking,       //                       .v_blanking
		output wire [15:0] avalon_camera_export_red_gain,         //                       .red_gain
		output wire [15:0] avalon_camera_export_blue_gain,        //                       .blue_gain
		output wire [15:0] avalon_camera_export_green1_gain,      //                       .green1_gain
		output wire [15:0] avalon_camera_export_green2_gain,      //                       .green2_gain
		input  wire        ccd_pixel_clock_bridge_clk,            // ccd_pixel_clock_bridge.clk
		input  wire        clk_50_clk,                            //                 clk_50.clk
		output wire        h2f_reset_reset_n,                     //              h2f_reset.reset_n
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK, //           hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,   //                       .hps_io_emac1_inst_TXD0
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,   //                       .hps_io_emac1_inst_TXD1
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,   //                       .hps_io_emac1_inst_TXD2
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,   //                       .hps_io_emac1_inst_TXD3
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,   //                       .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,   //                       .hps_io_emac1_inst_MDIO
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,    //                       .hps_io_emac1_inst_MDC
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL, //                       .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL, //                       .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK, //                       .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,   //                       .hps_io_emac1_inst_RXD1
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,   //                       .hps_io_emac1_inst_RXD2
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,   //                       .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,     //                       .hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,      //                       .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,      //                       .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,     //                       .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,      //                       .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,      //                       .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,      //                       .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,      //                       .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,      //                       .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,      //                       .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,      //                       .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,      //                       .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,      //                       .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,      //                       .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,     //                       .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,     //                       .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,     //                       .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,     //                       .hps_io_usb1_inst_NXT
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,     //                       .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,     //                       .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SDA,     //                       .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SCL,     //                       .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,  //                       .hps_io_gpio_inst_GPIO09
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,  //                       .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO40,  //                       .hps_io_gpio_inst_GPIO40
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,  //                       .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,  //                       .hps_io_gpio_inst_GPIO54
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO61,  //                       .hps_io_gpio_inst_GPIO61
		output wire [14:0] memory_mem_a,                          //                 memory.mem_a
		output wire [2:0]  memory_mem_ba,                         //                       .mem_ba
		output wire        memory_mem_ck,                         //                       .mem_ck
		output wire        memory_mem_ck_n,                       //                       .mem_ck_n
		output wire        memory_mem_cke,                        //                       .mem_cke
		output wire        memory_mem_cs_n,                       //                       .mem_cs_n
		output wire        memory_mem_ras_n,                      //                       .mem_ras_n
		output wire        memory_mem_cas_n,                      //                       .mem_cas_n
		output wire        memory_mem_we_n,                       //                       .mem_we_n
		output wire        memory_mem_reset_n,                    //                       .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                         //                       .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                        //                       .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                      //                       .mem_dqs_n
		output wire        memory_mem_odt,                        //                       .mem_odt
		output wire [3:0]  memory_mem_dm,                         //                       .mem_dm
		input  wire        memory_oct_rzqin,                      //                       .oct_rzqin
		output wire        pll_camera_clks_24_clk,                //     pll_camera_clks_24.clk
		output wire        pll_vga_clks_191_clk,                  //       pll_vga_clks_191.clk
		output wire        pll_vga_clks_25_clk,                   //        pll_vga_clks_25.clk
		input  wire        rgbgray_img_data_valid,                //            rgbgray_img.data_valid
		input  wire [31:0] rgbgray_img_input_data,                //                       .input_data
		input  wire [15:0] rgbgray_img_img_width,                 //                       .img_width
		input  wire [15:0] rgbgray_img_img_height,                //                       .img_height
		input  wire        rgbgray_stream_reset_n_reset_n         // rgbgray_stream_reset_n.reset_n
	);

	wire          hps_0_h2f_reset_reset;                                              // hps_0:h2f_rst_n -> [pll_camera_clks:rst, pll_vga_clks:rst, rst_controller:reset_in0]
	wire   [31:0] accel_0_avalon_master_readdata;                                     // mm_interconnect_0:accel_0_avalon_master_readdata -> accel_0:M_readdata
	wire          accel_0_avalon_master_waitrequest;                                  // mm_interconnect_0:accel_0_avalon_master_waitrequest -> accel_0:M_waitrequest
	wire   [31:0] accel_0_avalon_master_address;                                      // accel_0:M_address -> mm_interconnect_0:accel_0_avalon_master_address
	wire          accel_0_avalon_master_read;                                         // accel_0:M_read -> mm_interconnect_0:accel_0_avalon_master_read
	wire   [31:0] accel_0_avalon_master_writedata;                                    // accel_0:M_writedata -> mm_interconnect_0:accel_0_avalon_master_writedata
	wire          accel_0_avalon_master_write;                                        // accel_0:M_write -> mm_interconnect_0:accel_0_avalon_master_write
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_awburst;                      // mm_interconnect_0:hps_0_f2h_axi_slave_awburst -> hps_0:f2h_AWBURST
	wire    [4:0] mm_interconnect_0_hps_0_f2h_axi_slave_awuser;                       // mm_interconnect_0:hps_0_f2h_axi_slave_awuser -> hps_0:f2h_AWUSER
	wire    [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_arlen;                        // mm_interconnect_0:hps_0_f2h_axi_slave_arlen -> hps_0:f2h_ARLEN
	wire   [15:0] mm_interconnect_0_hps_0_f2h_axi_slave_wstrb;                        // mm_interconnect_0:hps_0_f2h_axi_slave_wstrb -> hps_0:f2h_WSTRB
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_wready;                       // hps_0:f2h_WREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_wready
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_rid;                          // hps_0:f2h_RID -> mm_interconnect_0:hps_0_f2h_axi_slave_rid
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_rready;                       // mm_interconnect_0:hps_0_f2h_axi_slave_rready -> hps_0:f2h_RREADY
	wire    [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_awlen;                        // mm_interconnect_0:hps_0_f2h_axi_slave_awlen -> hps_0:f2h_AWLEN
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_wid;                          // mm_interconnect_0:hps_0_f2h_axi_slave_wid -> hps_0:f2h_WID
	wire    [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_arcache;                      // mm_interconnect_0:hps_0_f2h_axi_slave_arcache -> hps_0:f2h_ARCACHE
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_wvalid;                       // mm_interconnect_0:hps_0_f2h_axi_slave_wvalid -> hps_0:f2h_WVALID
	wire   [31:0] mm_interconnect_0_hps_0_f2h_axi_slave_araddr;                       // mm_interconnect_0:hps_0_f2h_axi_slave_araddr -> hps_0:f2h_ARADDR
	wire    [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_arprot;                       // mm_interconnect_0:hps_0_f2h_axi_slave_arprot -> hps_0:f2h_ARPROT
	wire    [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_awprot;                       // mm_interconnect_0:hps_0_f2h_axi_slave_awprot -> hps_0:f2h_AWPROT
	wire  [127:0] mm_interconnect_0_hps_0_f2h_axi_slave_wdata;                        // mm_interconnect_0:hps_0_f2h_axi_slave_wdata -> hps_0:f2h_WDATA
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_arvalid;                      // mm_interconnect_0:hps_0_f2h_axi_slave_arvalid -> hps_0:f2h_ARVALID
	wire    [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_awcache;                      // mm_interconnect_0:hps_0_f2h_axi_slave_awcache -> hps_0:f2h_AWCACHE
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_arid;                         // mm_interconnect_0:hps_0_f2h_axi_slave_arid -> hps_0:f2h_ARID
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_arlock;                       // mm_interconnect_0:hps_0_f2h_axi_slave_arlock -> hps_0:f2h_ARLOCK
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_awlock;                       // mm_interconnect_0:hps_0_f2h_axi_slave_awlock -> hps_0:f2h_AWLOCK
	wire   [31:0] mm_interconnect_0_hps_0_f2h_axi_slave_awaddr;                       // mm_interconnect_0:hps_0_f2h_axi_slave_awaddr -> hps_0:f2h_AWADDR
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_bresp;                        // hps_0:f2h_BRESP -> mm_interconnect_0:hps_0_f2h_axi_slave_bresp
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_arready;                      // hps_0:f2h_ARREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_arready
	wire  [127:0] mm_interconnect_0_hps_0_f2h_axi_slave_rdata;                        // hps_0:f2h_RDATA -> mm_interconnect_0:hps_0_f2h_axi_slave_rdata
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_awready;                      // hps_0:f2h_AWREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_awready
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_arburst;                      // mm_interconnect_0:hps_0_f2h_axi_slave_arburst -> hps_0:f2h_ARBURST
	wire    [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_arsize;                       // mm_interconnect_0:hps_0_f2h_axi_slave_arsize -> hps_0:f2h_ARSIZE
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_bready;                       // mm_interconnect_0:hps_0_f2h_axi_slave_bready -> hps_0:f2h_BREADY
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_rlast;                        // hps_0:f2h_RLAST -> mm_interconnect_0:hps_0_f2h_axi_slave_rlast
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_wlast;                        // mm_interconnect_0:hps_0_f2h_axi_slave_wlast -> hps_0:f2h_WLAST
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_rresp;                        // hps_0:f2h_RRESP -> mm_interconnect_0:hps_0_f2h_axi_slave_rresp
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_awid;                         // mm_interconnect_0:hps_0_f2h_axi_slave_awid -> hps_0:f2h_AWID
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_bid;                          // hps_0:f2h_BID -> mm_interconnect_0:hps_0_f2h_axi_slave_bid
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_bvalid;                       // hps_0:f2h_BVALID -> mm_interconnect_0:hps_0_f2h_axi_slave_bvalid
	wire    [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_awsize;                       // mm_interconnect_0:hps_0_f2h_axi_slave_awsize -> hps_0:f2h_AWSIZE
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_awvalid;                      // mm_interconnect_0:hps_0_f2h_axi_slave_awvalid -> hps_0:f2h_AWVALID
	wire    [4:0] mm_interconnect_0_hps_0_f2h_axi_slave_aruser;                       // mm_interconnect_0:hps_0_f2h_axi_slave_aruser -> hps_0:f2h_ARUSER
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_rvalid;                       // hps_0:f2h_RVALID -> mm_interconnect_0:hps_0_f2h_axi_slave_rvalid
	wire          avalon_img_writer_rgbgray_avalon_master_waitrequest;                // mm_interconnect_1:avalon_img_writer_rgbgray_avalon_master_waitrequest -> avalon_img_writer_rgbgray:M_waitrequest
	wire   [31:0] avalon_img_writer_rgbgray_avalon_master_address;                    // avalon_img_writer_rgbgray:M_address -> mm_interconnect_1:avalon_img_writer_rgbgray_avalon_master_address
	wire   [15:0] avalon_img_writer_rgbgray_avalon_master_byteenable;                 // avalon_img_writer_rgbgray:M_byteenable -> mm_interconnect_1:avalon_img_writer_rgbgray_avalon_master_byteenable
	wire          avalon_img_writer_rgbgray_avalon_master_write;                      // avalon_img_writer_rgbgray:M_write -> mm_interconnect_1:avalon_img_writer_rgbgray_avalon_master_write
	wire  [127:0] avalon_img_writer_rgbgray_avalon_master_writedata;                  // avalon_img_writer_rgbgray:M_writedata -> mm_interconnect_1:avalon_img_writer_rgbgray_avalon_master_writedata
	wire    [6:0] avalon_img_writer_rgbgray_avalon_master_burstcount;                 // avalon_img_writer_rgbgray:M_burstcount -> mm_interconnect_1:avalon_img_writer_rgbgray_avalon_master_burstcount
	wire          mm_interconnect_1_hps_0_f2h_sdram1_data_waitrequest;                // hps_0:f2h_sdram1_WAITREQUEST -> mm_interconnect_1:hps_0_f2h_sdram1_data_waitrequest
	wire   [27:0] mm_interconnect_1_hps_0_f2h_sdram1_data_address;                    // mm_interconnect_1:hps_0_f2h_sdram1_data_address -> hps_0:f2h_sdram1_ADDRESS
	wire   [15:0] mm_interconnect_1_hps_0_f2h_sdram1_data_byteenable;                 // mm_interconnect_1:hps_0_f2h_sdram1_data_byteenable -> hps_0:f2h_sdram1_BYTEENABLE
	wire          mm_interconnect_1_hps_0_f2h_sdram1_data_write;                      // mm_interconnect_1:hps_0_f2h_sdram1_data_write -> hps_0:f2h_sdram1_WRITE
	wire  [127:0] mm_interconnect_1_hps_0_f2h_sdram1_data_writedata;                  // mm_interconnect_1:hps_0_f2h_sdram1_data_writedata -> hps_0:f2h_sdram1_WRITEDATA
	wire    [7:0] mm_interconnect_1_hps_0_f2h_sdram1_data_burstcount;                 // mm_interconnect_1:hps_0_f2h_sdram1_data_burstcount -> hps_0:f2h_sdram1_BURSTCOUNT
	wire    [1:0] hps_0_h2f_axi_master_awburst;                                       // hps_0:h2f_AWBURST -> mm_interconnect_2:hps_0_h2f_axi_master_awburst
	wire    [3:0] hps_0_h2f_axi_master_arlen;                                         // hps_0:h2f_ARLEN -> mm_interconnect_2:hps_0_h2f_axi_master_arlen
	wire   [15:0] hps_0_h2f_axi_master_wstrb;                                         // hps_0:h2f_WSTRB -> mm_interconnect_2:hps_0_h2f_axi_master_wstrb
	wire          hps_0_h2f_axi_master_wready;                                        // mm_interconnect_2:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire   [11:0] hps_0_h2f_axi_master_rid;                                           // mm_interconnect_2:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_rready;                                        // hps_0:h2f_RREADY -> mm_interconnect_2:hps_0_h2f_axi_master_rready
	wire    [3:0] hps_0_h2f_axi_master_awlen;                                         // hps_0:h2f_AWLEN -> mm_interconnect_2:hps_0_h2f_axi_master_awlen
	wire   [11:0] hps_0_h2f_axi_master_wid;                                           // hps_0:h2f_WID -> mm_interconnect_2:hps_0_h2f_axi_master_wid
	wire    [3:0] hps_0_h2f_axi_master_arcache;                                       // hps_0:h2f_ARCACHE -> mm_interconnect_2:hps_0_h2f_axi_master_arcache
	wire          hps_0_h2f_axi_master_wvalid;                                        // hps_0:h2f_WVALID -> mm_interconnect_2:hps_0_h2f_axi_master_wvalid
	wire   [29:0] hps_0_h2f_axi_master_araddr;                                        // hps_0:h2f_ARADDR -> mm_interconnect_2:hps_0_h2f_axi_master_araddr
	wire    [2:0] hps_0_h2f_axi_master_arprot;                                        // hps_0:h2f_ARPROT -> mm_interconnect_2:hps_0_h2f_axi_master_arprot
	wire    [2:0] hps_0_h2f_axi_master_awprot;                                        // hps_0:h2f_AWPROT -> mm_interconnect_2:hps_0_h2f_axi_master_awprot
	wire  [127:0] hps_0_h2f_axi_master_wdata;                                         // hps_0:h2f_WDATA -> mm_interconnect_2:hps_0_h2f_axi_master_wdata
	wire          hps_0_h2f_axi_master_arvalid;                                       // hps_0:h2f_ARVALID -> mm_interconnect_2:hps_0_h2f_axi_master_arvalid
	wire    [3:0] hps_0_h2f_axi_master_awcache;                                       // hps_0:h2f_AWCACHE -> mm_interconnect_2:hps_0_h2f_axi_master_awcache
	wire   [11:0] hps_0_h2f_axi_master_arid;                                          // hps_0:h2f_ARID -> mm_interconnect_2:hps_0_h2f_axi_master_arid
	wire    [1:0] hps_0_h2f_axi_master_arlock;                                        // hps_0:h2f_ARLOCK -> mm_interconnect_2:hps_0_h2f_axi_master_arlock
	wire    [1:0] hps_0_h2f_axi_master_awlock;                                        // hps_0:h2f_AWLOCK -> mm_interconnect_2:hps_0_h2f_axi_master_awlock
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                                        // hps_0:h2f_AWADDR -> mm_interconnect_2:hps_0_h2f_axi_master_awaddr
	wire    [1:0] hps_0_h2f_axi_master_bresp;                                         // mm_interconnect_2:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire          hps_0_h2f_axi_master_arready;                                       // mm_interconnect_2:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [127:0] hps_0_h2f_axi_master_rdata;                                         // mm_interconnect_2:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire          hps_0_h2f_axi_master_awready;                                       // mm_interconnect_2:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                                       // hps_0:h2f_ARBURST -> mm_interconnect_2:hps_0_h2f_axi_master_arburst
	wire    [2:0] hps_0_h2f_axi_master_arsize;                                        // hps_0:h2f_ARSIZE -> mm_interconnect_2:hps_0_h2f_axi_master_arsize
	wire          hps_0_h2f_axi_master_bready;                                        // hps_0:h2f_BREADY -> mm_interconnect_2:hps_0_h2f_axi_master_bready
	wire          hps_0_h2f_axi_master_rlast;                                         // mm_interconnect_2:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire          hps_0_h2f_axi_master_wlast;                                         // hps_0:h2f_WLAST -> mm_interconnect_2:hps_0_h2f_axi_master_wlast
	wire    [1:0] hps_0_h2f_axi_master_rresp;                                         // mm_interconnect_2:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire   [11:0] hps_0_h2f_axi_master_awid;                                          // hps_0:h2f_AWID -> mm_interconnect_2:hps_0_h2f_axi_master_awid
	wire   [11:0] hps_0_h2f_axi_master_bid;                                           // mm_interconnect_2:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire          hps_0_h2f_axi_master_bvalid;                                        // mm_interconnect_2:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire    [2:0] hps_0_h2f_axi_master_awsize;                                        // hps_0:h2f_AWSIZE -> mm_interconnect_2:hps_0_h2f_axi_master_awsize
	wire          hps_0_h2f_axi_master_awvalid;                                       // hps_0:h2f_AWVALID -> mm_interconnect_2:hps_0_h2f_axi_master_awvalid
	wire          hps_0_h2f_axi_master_rvalid;                                        // mm_interconnect_2:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire   [31:0] mm_interconnect_2_avalon_img_writer_rgbgray_avalon_slave_readdata;  // avalon_img_writer_rgbgray:S_readdata -> mm_interconnect_2:avalon_img_writer_rgbgray_avalon_slave_readdata
	wire    [3:0] mm_interconnect_2_avalon_img_writer_rgbgray_avalon_slave_address;   // mm_interconnect_2:avalon_img_writer_rgbgray_avalon_slave_address -> avalon_img_writer_rgbgray:S_address
	wire          mm_interconnect_2_avalon_img_writer_rgbgray_avalon_slave_read;      // mm_interconnect_2:avalon_img_writer_rgbgray_avalon_slave_read -> avalon_img_writer_rgbgray:S_read
	wire          mm_interconnect_2_avalon_img_writer_rgbgray_avalon_slave_write;     // mm_interconnect_2:avalon_img_writer_rgbgray_avalon_slave_write -> avalon_img_writer_rgbgray:S_write
	wire   [31:0] mm_interconnect_2_avalon_img_writer_rgbgray_avalon_slave_writedata; // mm_interconnect_2:avalon_img_writer_rgbgray_avalon_slave_writedata -> avalon_img_writer_rgbgray:S_writedata
	wire   [31:0] mm_interconnect_2_accel_0_avalon_slave_readdata;                    // accel_0:S_readdata -> mm_interconnect_2:accel_0_avalon_slave_readdata
	wire          mm_interconnect_2_accel_0_avalon_slave_waitrequest;                 // accel_0:S_waitrequest -> mm_interconnect_2:accel_0_avalon_slave_waitrequest
	wire    [2:0] mm_interconnect_2_accel_0_avalon_slave_address;                     // mm_interconnect_2:accel_0_avalon_slave_address -> accel_0:S_address
	wire          mm_interconnect_2_accel_0_avalon_slave_read;                        // mm_interconnect_2:accel_0_avalon_slave_read -> accel_0:S_read
	wire          mm_interconnect_2_accel_0_avalon_slave_write;                       // mm_interconnect_2:accel_0_avalon_slave_write -> accel_0:S_write
	wire   [31:0] mm_interconnect_2_accel_0_avalon_slave_writedata;                   // mm_interconnect_2:accel_0_avalon_slave_writedata -> accel_0:S_writedata
	wire   [31:0] mm_interconnect_2_avalon_camera_0_s1_readdata;                      // avalon_camera_0:avs_s1_readdata -> mm_interconnect_2:avalon_camera_0_s1_readdata
	wire    [4:0] mm_interconnect_2_avalon_camera_0_s1_address;                       // mm_interconnect_2:avalon_camera_0_s1_address -> avalon_camera_0:avs_s1_address
	wire          mm_interconnect_2_avalon_camera_0_s1_read;                          // mm_interconnect_2:avalon_camera_0_s1_read -> avalon_camera_0:avs_s1_read
	wire          mm_interconnect_2_avalon_camera_0_s1_write;                         // mm_interconnect_2:avalon_camera_0_s1_write -> avalon_camera_0:avs_s1_write
	wire   [31:0] mm_interconnect_2_avalon_camera_0_s1_writedata;                     // mm_interconnect_2:avalon_camera_0_s1_writedata -> avalon_camera_0:avs_s1_writedata
	wire   [31:0] hps_0_f2h_irq0_irq;                                                 // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                                 // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire          rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [accel_0:rst_n, avalon_camera_0:reset_n, avalon_img_writer_rgbgray:reset_n, mm_interconnect_0:accel_0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:avalon_img_writer_rgbgray_reset_reset_bridge_in_reset_reset, mm_interconnect_2:avalon_img_writer_rgbgray_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]

	accel accel_0 (
		.clk           (ccd_pixel_clock_bridge_clk),                         //         clock.clk
		.M_address     (accel_0_avalon_master_address),                      // avalon_master.address
		.M_writedata   (accel_0_avalon_master_writedata),                    //              .writedata
		.M_write       (accel_0_avalon_master_write),                        //              .write
		.M_readdata    (accel_0_avalon_master_readdata),                     //              .readdata
		.M_read        (accel_0_avalon_master_read),                         //              .read
		.M_waitrequest (accel_0_avalon_master_waitrequest),                  //              .waitrequest
		.rst_n         (~rst_controller_reset_out_reset),                    //    reset_sink.reset_n
		.S_address     (mm_interconnect_2_accel_0_avalon_slave_address),     //  avalon_slave.address
		.S_writedata   (mm_interconnect_2_accel_0_avalon_slave_writedata),   //              .writedata
		.S_write       (mm_interconnect_2_accel_0_avalon_slave_write),       //              .write
		.S_readdata    (mm_interconnect_2_accel_0_avalon_slave_readdata),    //              .readdata
		.S_read        (mm_interconnect_2_accel_0_avalon_slave_read),        //              .read
		.S_waitrequest (mm_interconnect_2_accel_0_avalon_slave_waitrequest)  //              .waitrequest
	);

	avalon_camera #(
		.WIDTH        (18'b000000001010000000),
		.HEIGHT       (18'b000000000111100000),
		.START_ROW    (18'b000000000000000000),
		.START_COLUMN (18'b000000000000000000),
		.ROW_SIZE     (18'b000000011101111111),
		.COLUMN_SIZE  (18'b000000100111111111),
		.ROW_MODE     (18'b000000000000000011),
		.COLUMN_MODE  (18'b000000000000000011),
		.EXPOSURE     (18'b000000001111111111),
		.H_BLANKING   (18'b000000000000000000),
		.V_BLANKING   (18'b000000000000011001),
		.RED_GAIN     (18'b000000000010011100),
		.BLUE_GAIN    (18'b000000000010011010),
		.GREEN1_GAIN  (18'b000000000000010011),
		.GREEN2_GAIN  (18'b000000000000010011)
	) avalon_camera_0 (
		.clk                         (ccd_pixel_clock_bridge_clk),                     //  clock.clk
		.avs_export_height           (avalon_camera_export_height),                    // export.height
		.avs_export_start_row        (avalon_camera_export_startrow),                  //       .startrow
		.avs_export_start_column     (avalon_camera_export_startcol),                  //       .startcol
		.avs_export_column_mode      (avalon_camera_export_colmode),                   //       .colmode
		.avs_export_exposure         (avalon_camera_export_exposure),                  //       .exposure
		.avs_export_row_size         (avalon_camera_export_rowsize),                   //       .rowsize
		.avs_export_column_size      (avalon_camera_export_colsize),                   //       .colsize
		.avs_export_row_mode         (avalon_camera_export_rowmode),                   //       .rowmode
		.avs_export_cam_soft_reset_n (avalon_camera_export_soft_reset_n),              //       .soft_reset_n
		.avs_export_width            (avalon_camera_export_width),                     //       .width
		.avs_export_h_blanking       (avalon_camera_export_h_blanking),                //       .h_blanking
		.avs_export_v_blanking       (avalon_camera_export_v_blanking),                //       .v_blanking
		.avs_export_red_gain         (avalon_camera_export_red_gain),                  //       .red_gain
		.avs_export_blue_gain        (avalon_camera_export_blue_gain),                 //       .blue_gain
		.avs_export_green1_gain      (avalon_camera_export_green1_gain),               //       .green1_gain
		.avs_export_green2_gain      (avalon_camera_export_green2_gain),               //       .green2_gain
		.reset_n                     (~rst_controller_reset_out_reset),                //  reset.reset_n
		.avs_s1_address              (mm_interconnect_2_avalon_camera_0_s1_address),   //     s1.address
		.avs_s1_read                 (mm_interconnect_2_avalon_camera_0_s1_read),      //       .read
		.avs_s1_readdata             (mm_interconnect_2_avalon_camera_0_s1_readdata),  //       .readdata
		.avs_s1_write                (mm_interconnect_2_avalon_camera_0_s1_write),     //       .write
		.avs_s1_writedata            (mm_interconnect_2_avalon_camera_0_s1_writedata)  //       .writedata
	);

	avalon_image_writer #(
		.COMPONENT_SIZE    (8),
		.NUMBER_COMPONENTS (4),
		.PIX_WR            (4)
	) avalon_img_writer_rgbgray (
		.clk            (ccd_pixel_clock_bridge_clk),                                         //             clock.clk
		.reset_n        (~rst_controller_reset_out_reset),                                    //             reset.reset_n
		.S_address      (mm_interconnect_2_avalon_img_writer_rgbgray_avalon_slave_address),   //      avalon_slave.address
		.S_writedata    (mm_interconnect_2_avalon_img_writer_rgbgray_avalon_slave_writedata), //                  .writedata
		.S_readdata     (mm_interconnect_2_avalon_img_writer_rgbgray_avalon_slave_readdata),  //                  .readdata
		.S_write        (mm_interconnect_2_avalon_img_writer_rgbgray_avalon_slave_write),     //                  .write
		.S_read         (mm_interconnect_2_avalon_img_writer_rgbgray_avalon_slave_read),      //                  .read
		.M_address      (avalon_img_writer_rgbgray_avalon_master_address),                    //     avalon_master.address
		.M_write        (avalon_img_writer_rgbgray_avalon_master_write),                      //                  .write
		.M_byteenable   (avalon_img_writer_rgbgray_avalon_master_byteenable),                 //                  .byteenable
		.M_writedata    (avalon_img_writer_rgbgray_avalon_master_writedata),                  //                  .writedata
		.M_waitrequest  (avalon_img_writer_rgbgray_avalon_master_waitrequest),                //                  .waitrequest
		.M_burstcount   (avalon_img_writer_rgbgray_avalon_master_burstcount),                 //                  .burstcount
		.data_valid     (rgbgray_img_data_valid),                                             //       conduit_end.data_valid
		.input_data     (rgbgray_img_input_data),                                             //                  .input_data
		.img_width      (rgbgray_img_img_width),                                              //                  .img_width
		.img_height     (rgbgray_img_img_height),                                             //                  .img_height
		.stream_reset_n (rgbgray_stream_reset_n_reset_n)                                      // stream_reset_sink.reset_n
	);

	soc_system_hps_0 #(
		.F2S_Width (3),
		.S2F_Width (3)
	) hps_0 (
		.mem_a                    (memory_mem_a),                                        //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                                       //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                                       //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                                     //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                      //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                                     //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                                    //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                                    //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                                     //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                                  //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                       //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                      //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                                    //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                      //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                                       //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                                    //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_0_hps_io_hps_io_emac1_inst_TX_CLK),               //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_0_hps_io_hps_io_emac1_inst_TXD0),                 //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_0_hps_io_hps_io_emac1_inst_TXD1),                 //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_0_hps_io_hps_io_emac1_inst_TXD2),                 //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_0_hps_io_hps_io_emac1_inst_TXD3),                 //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_0_hps_io_hps_io_emac1_inst_RXD0),                 //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_0_hps_io_hps_io_emac1_inst_MDIO),                 //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_0_hps_io_hps_io_emac1_inst_MDC),                  //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_0_hps_io_hps_io_emac1_inst_RX_CTL),               //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_0_hps_io_hps_io_emac1_inst_TX_CTL),               //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_0_hps_io_hps_io_emac1_inst_RX_CLK),               //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_0_hps_io_hps_io_emac1_inst_RXD1),                 //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_0_hps_io_hps_io_emac1_inst_RXD2),                 //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_0_hps_io_hps_io_emac1_inst_RXD3),                 //                  .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_0_hps_io_hps_io_sdio_inst_CMD),                   //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_0_hps_io_hps_io_sdio_inst_D0),                    //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_0_hps_io_hps_io_sdio_inst_D1),                    //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_0_hps_io_hps_io_sdio_inst_CLK),                   //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_0_hps_io_hps_io_sdio_inst_D2),                    //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_0_hps_io_hps_io_sdio_inst_D3),                    //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_0_hps_io_hps_io_usb1_inst_D0),                    //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_0_hps_io_hps_io_usb1_inst_D1),                    //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_0_hps_io_hps_io_usb1_inst_D2),                    //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_0_hps_io_hps_io_usb1_inst_D3),                    //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_0_hps_io_hps_io_usb1_inst_D4),                    //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_0_hps_io_hps_io_usb1_inst_D5),                    //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_0_hps_io_hps_io_usb1_inst_D6),                    //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_0_hps_io_hps_io_usb1_inst_D7),                    //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_0_hps_io_hps_io_usb1_inst_CLK),                   //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_0_hps_io_hps_io_usb1_inst_STP),                   //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_0_hps_io_hps_io_usb1_inst_DIR),                   //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_0_hps_io_hps_io_usb1_inst_NXT),                   //                  .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX     (hps_0_hps_io_hps_io_uart0_inst_RX),                   //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_0_hps_io_hps_io_uart0_inst_TX),                   //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_0_hps_io_hps_io_i2c0_inst_SDA),                   //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_0_hps_io_hps_io_i2c0_inst_SCL),                   //                  .hps_io_i2c0_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_0_hps_io_hps_io_gpio_inst_GPIO09),                //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_0_hps_io_hps_io_gpio_inst_GPIO35),                //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_0_hps_io_hps_io_gpio_inst_GPIO40),                //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO53  (hps_0_hps_io_hps_io_gpio_inst_GPIO53),                //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_0_hps_io_hps_io_gpio_inst_GPIO54),                //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_0_hps_io_hps_io_gpio_inst_GPIO61),                //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset),                               //         h2f_reset.reset_n
		.f2h_sdram0_clk           (ccd_pixel_clock_bridge_clk),                          //  f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (),                                                    //   f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (),                                                    //                  .burstcount
		.f2h_sdram0_WAITREQUEST   (),                                                    //                  .waitrequest
		.f2h_sdram0_READDATA      (),                                                    //                  .readdata
		.f2h_sdram0_READDATAVALID (),                                                    //                  .readdatavalid
		.f2h_sdram0_READ          (),                                                    //                  .read
		.f2h_sdram0_WRITEDATA     (),                                                    //                  .writedata
		.f2h_sdram0_BYTEENABLE    (),                                                    //                  .byteenable
		.f2h_sdram0_WRITE         (),                                                    //                  .write
		.f2h_sdram1_clk           (ccd_pixel_clock_bridge_clk),                          //  f2h_sdram1_clock.clk
		.f2h_sdram1_ADDRESS       (mm_interconnect_1_hps_0_f2h_sdram1_data_address),     //   f2h_sdram1_data.address
		.f2h_sdram1_BURSTCOUNT    (mm_interconnect_1_hps_0_f2h_sdram1_data_burstcount),  //                  .burstcount
		.f2h_sdram1_WAITREQUEST   (mm_interconnect_1_hps_0_f2h_sdram1_data_waitrequest), //                  .waitrequest
		.f2h_sdram1_WRITEDATA     (mm_interconnect_1_hps_0_f2h_sdram1_data_writedata),   //                  .writedata
		.f2h_sdram1_BYTEENABLE    (mm_interconnect_1_hps_0_f2h_sdram1_data_byteenable),  //                  .byteenable
		.f2h_sdram1_WRITE         (mm_interconnect_1_hps_0_f2h_sdram1_data_write),       //                  .write
		.h2f_axi_clk              (ccd_pixel_clock_bridge_clk),                          //     h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),                           //    h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),                         //                  .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),                          //                  .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),                         //                  .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),                        //                  .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),                         //                  .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),                        //                  .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),                         //                  .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),                        //                  .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),                        //                  .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),                            //                  .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),                          //                  .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),                          //                  .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),                          //                  .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),                         //                  .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),                         //                  .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),                            //                  .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),                          //                  .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),                         //                  .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),                         //                  .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),                           //                  .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),                         //                  .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),                          //                  .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),                         //                  .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),                        //                  .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),                         //                  .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),                        //                  .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),                         //                  .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),                        //                  .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),                        //                  .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),                            //                  .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),                          //                  .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),                          //                  .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),                          //                  .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),                         //                  .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready),                         //                  .rready
		.f2h_axi_clk              (ccd_pixel_clock_bridge_clk),                          //     f2h_axi_clock.clk
		.f2h_AWID                 (mm_interconnect_0_hps_0_f2h_axi_slave_awid),          //     f2h_axi_slave.awid
		.f2h_AWADDR               (mm_interconnect_0_hps_0_f2h_axi_slave_awaddr),        //                  .awaddr
		.f2h_AWLEN                (mm_interconnect_0_hps_0_f2h_axi_slave_awlen),         //                  .awlen
		.f2h_AWSIZE               (mm_interconnect_0_hps_0_f2h_axi_slave_awsize),        //                  .awsize
		.f2h_AWBURST              (mm_interconnect_0_hps_0_f2h_axi_slave_awburst),       //                  .awburst
		.f2h_AWLOCK               (mm_interconnect_0_hps_0_f2h_axi_slave_awlock),        //                  .awlock
		.f2h_AWCACHE              (mm_interconnect_0_hps_0_f2h_axi_slave_awcache),       //                  .awcache
		.f2h_AWPROT               (mm_interconnect_0_hps_0_f2h_axi_slave_awprot),        //                  .awprot
		.f2h_AWVALID              (mm_interconnect_0_hps_0_f2h_axi_slave_awvalid),       //                  .awvalid
		.f2h_AWREADY              (mm_interconnect_0_hps_0_f2h_axi_slave_awready),       //                  .awready
		.f2h_AWUSER               (mm_interconnect_0_hps_0_f2h_axi_slave_awuser),        //                  .awuser
		.f2h_WID                  (mm_interconnect_0_hps_0_f2h_axi_slave_wid),           //                  .wid
		.f2h_WDATA                (mm_interconnect_0_hps_0_f2h_axi_slave_wdata),         //                  .wdata
		.f2h_WSTRB                (mm_interconnect_0_hps_0_f2h_axi_slave_wstrb),         //                  .wstrb
		.f2h_WLAST                (mm_interconnect_0_hps_0_f2h_axi_slave_wlast),         //                  .wlast
		.f2h_WVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_wvalid),        //                  .wvalid
		.f2h_WREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_wready),        //                  .wready
		.f2h_BID                  (mm_interconnect_0_hps_0_f2h_axi_slave_bid),           //                  .bid
		.f2h_BRESP                (mm_interconnect_0_hps_0_f2h_axi_slave_bresp),         //                  .bresp
		.f2h_BVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_bvalid),        //                  .bvalid
		.f2h_BREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_bready),        //                  .bready
		.f2h_ARID                 (mm_interconnect_0_hps_0_f2h_axi_slave_arid),          //                  .arid
		.f2h_ARADDR               (mm_interconnect_0_hps_0_f2h_axi_slave_araddr),        //                  .araddr
		.f2h_ARLEN                (mm_interconnect_0_hps_0_f2h_axi_slave_arlen),         //                  .arlen
		.f2h_ARSIZE               (mm_interconnect_0_hps_0_f2h_axi_slave_arsize),        //                  .arsize
		.f2h_ARBURST              (mm_interconnect_0_hps_0_f2h_axi_slave_arburst),       //                  .arburst
		.f2h_ARLOCK               (mm_interconnect_0_hps_0_f2h_axi_slave_arlock),        //                  .arlock
		.f2h_ARCACHE              (mm_interconnect_0_hps_0_f2h_axi_slave_arcache),       //                  .arcache
		.f2h_ARPROT               (mm_interconnect_0_hps_0_f2h_axi_slave_arprot),        //                  .arprot
		.f2h_ARVALID              (mm_interconnect_0_hps_0_f2h_axi_slave_arvalid),       //                  .arvalid
		.f2h_ARREADY              (mm_interconnect_0_hps_0_f2h_axi_slave_arready),       //                  .arready
		.f2h_ARUSER               (mm_interconnect_0_hps_0_f2h_axi_slave_aruser),        //                  .aruser
		.f2h_RID                  (mm_interconnect_0_hps_0_f2h_axi_slave_rid),           //                  .rid
		.f2h_RDATA                (mm_interconnect_0_hps_0_f2h_axi_slave_rdata),         //                  .rdata
		.f2h_RRESP                (mm_interconnect_0_hps_0_f2h_axi_slave_rresp),         //                  .rresp
		.f2h_RLAST                (mm_interconnect_0_hps_0_f2h_axi_slave_rlast),         //                  .rlast
		.f2h_RVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_rvalid),        //                  .rvalid
		.f2h_RREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_rready),        //                  .rready
		.h2f_lw_axi_clk           (ccd_pixel_clock_bridge_clk),                          //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (),                                                    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (),                                                    //                  .awaddr
		.h2f_lw_AWLEN             (),                                                    //                  .awlen
		.h2f_lw_AWSIZE            (),                                                    //                  .awsize
		.h2f_lw_AWBURST           (),                                                    //                  .awburst
		.h2f_lw_AWLOCK            (),                                                    //                  .awlock
		.h2f_lw_AWCACHE           (),                                                    //                  .awcache
		.h2f_lw_AWPROT            (),                                                    //                  .awprot
		.h2f_lw_AWVALID           (),                                                    //                  .awvalid
		.h2f_lw_AWREADY           (),                                                    //                  .awready
		.h2f_lw_WID               (),                                                    //                  .wid
		.h2f_lw_WDATA             (),                                                    //                  .wdata
		.h2f_lw_WSTRB             (),                                                    //                  .wstrb
		.h2f_lw_WLAST             (),                                                    //                  .wlast
		.h2f_lw_WVALID            (),                                                    //                  .wvalid
		.h2f_lw_WREADY            (),                                                    //                  .wready
		.h2f_lw_BID               (),                                                    //                  .bid
		.h2f_lw_BRESP             (),                                                    //                  .bresp
		.h2f_lw_BVALID            (),                                                    //                  .bvalid
		.h2f_lw_BREADY            (),                                                    //                  .bready
		.h2f_lw_ARID              (),                                                    //                  .arid
		.h2f_lw_ARADDR            (),                                                    //                  .araddr
		.h2f_lw_ARLEN             (),                                                    //                  .arlen
		.h2f_lw_ARSIZE            (),                                                    //                  .arsize
		.h2f_lw_ARBURST           (),                                                    //                  .arburst
		.h2f_lw_ARLOCK            (),                                                    //                  .arlock
		.h2f_lw_ARCACHE           (),                                                    //                  .arcache
		.h2f_lw_ARPROT            (),                                                    //                  .arprot
		.h2f_lw_ARVALID           (),                                                    //                  .arvalid
		.h2f_lw_ARREADY           (),                                                    //                  .arready
		.h2f_lw_RID               (),                                                    //                  .rid
		.h2f_lw_RDATA             (),                                                    //                  .rdata
		.h2f_lw_RRESP             (),                                                    //                  .rresp
		.h2f_lw_RLAST             (),                                                    //                  .rlast
		.h2f_lw_RVALID            (),                                                    //                  .rvalid
		.h2f_lw_RREADY            (),                                                    //                  .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                                  //          f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                                   //          f2h_irq1.irq
	);

	soc_system_pll_camera_clks pll_camera_clks (
		.refclk   (clk_50_clk),             //  refclk.clk
		.rst      (~hps_0_h2f_reset_reset), //   reset.reset
		.outclk_0 (pll_camera_clks_24_clk), // outclk0.clk
		.locked   ()                        // (terminated)
	);

	soc_system_pll_vga_clks pll_vga_clks (
		.refclk   (clk_50_clk),             //  refclk.clk
		.rst      (~hps_0_h2f_reset_reset), //   reset.reset
		.outclk_0 (pll_vga_clks_25_clk),    // outclk0.clk
		.outclk_1 (pll_vga_clks_191_clk),   // outclk1.clk
		.locked   ()                        // (terminated)
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_f2h_axi_slave_awid                       (mm_interconnect_0_hps_0_f2h_axi_slave_awid),    //                      hps_0_f2h_axi_slave.awid
		.hps_0_f2h_axi_slave_awaddr                     (mm_interconnect_0_hps_0_f2h_axi_slave_awaddr),  //                                         .awaddr
		.hps_0_f2h_axi_slave_awlen                      (mm_interconnect_0_hps_0_f2h_axi_slave_awlen),   //                                         .awlen
		.hps_0_f2h_axi_slave_awsize                     (mm_interconnect_0_hps_0_f2h_axi_slave_awsize),  //                                         .awsize
		.hps_0_f2h_axi_slave_awburst                    (mm_interconnect_0_hps_0_f2h_axi_slave_awburst), //                                         .awburst
		.hps_0_f2h_axi_slave_awlock                     (mm_interconnect_0_hps_0_f2h_axi_slave_awlock),  //                                         .awlock
		.hps_0_f2h_axi_slave_awcache                    (mm_interconnect_0_hps_0_f2h_axi_slave_awcache), //                                         .awcache
		.hps_0_f2h_axi_slave_awprot                     (mm_interconnect_0_hps_0_f2h_axi_slave_awprot),  //                                         .awprot
		.hps_0_f2h_axi_slave_awuser                     (mm_interconnect_0_hps_0_f2h_axi_slave_awuser),  //                                         .awuser
		.hps_0_f2h_axi_slave_awvalid                    (mm_interconnect_0_hps_0_f2h_axi_slave_awvalid), //                                         .awvalid
		.hps_0_f2h_axi_slave_awready                    (mm_interconnect_0_hps_0_f2h_axi_slave_awready), //                                         .awready
		.hps_0_f2h_axi_slave_wid                        (mm_interconnect_0_hps_0_f2h_axi_slave_wid),     //                                         .wid
		.hps_0_f2h_axi_slave_wdata                      (mm_interconnect_0_hps_0_f2h_axi_slave_wdata),   //                                         .wdata
		.hps_0_f2h_axi_slave_wstrb                      (mm_interconnect_0_hps_0_f2h_axi_slave_wstrb),   //                                         .wstrb
		.hps_0_f2h_axi_slave_wlast                      (mm_interconnect_0_hps_0_f2h_axi_slave_wlast),   //                                         .wlast
		.hps_0_f2h_axi_slave_wvalid                     (mm_interconnect_0_hps_0_f2h_axi_slave_wvalid),  //                                         .wvalid
		.hps_0_f2h_axi_slave_wready                     (mm_interconnect_0_hps_0_f2h_axi_slave_wready),  //                                         .wready
		.hps_0_f2h_axi_slave_bid                        (mm_interconnect_0_hps_0_f2h_axi_slave_bid),     //                                         .bid
		.hps_0_f2h_axi_slave_bresp                      (mm_interconnect_0_hps_0_f2h_axi_slave_bresp),   //                                         .bresp
		.hps_0_f2h_axi_slave_bvalid                     (mm_interconnect_0_hps_0_f2h_axi_slave_bvalid),  //                                         .bvalid
		.hps_0_f2h_axi_slave_bready                     (mm_interconnect_0_hps_0_f2h_axi_slave_bready),  //                                         .bready
		.hps_0_f2h_axi_slave_arid                       (mm_interconnect_0_hps_0_f2h_axi_slave_arid),    //                                         .arid
		.hps_0_f2h_axi_slave_araddr                     (mm_interconnect_0_hps_0_f2h_axi_slave_araddr),  //                                         .araddr
		.hps_0_f2h_axi_slave_arlen                      (mm_interconnect_0_hps_0_f2h_axi_slave_arlen),   //                                         .arlen
		.hps_0_f2h_axi_slave_arsize                     (mm_interconnect_0_hps_0_f2h_axi_slave_arsize),  //                                         .arsize
		.hps_0_f2h_axi_slave_arburst                    (mm_interconnect_0_hps_0_f2h_axi_slave_arburst), //                                         .arburst
		.hps_0_f2h_axi_slave_arlock                     (mm_interconnect_0_hps_0_f2h_axi_slave_arlock),  //                                         .arlock
		.hps_0_f2h_axi_slave_arcache                    (mm_interconnect_0_hps_0_f2h_axi_slave_arcache), //                                         .arcache
		.hps_0_f2h_axi_slave_arprot                     (mm_interconnect_0_hps_0_f2h_axi_slave_arprot),  //                                         .arprot
		.hps_0_f2h_axi_slave_aruser                     (mm_interconnect_0_hps_0_f2h_axi_slave_aruser),  //                                         .aruser
		.hps_0_f2h_axi_slave_arvalid                    (mm_interconnect_0_hps_0_f2h_axi_slave_arvalid), //                                         .arvalid
		.hps_0_f2h_axi_slave_arready                    (mm_interconnect_0_hps_0_f2h_axi_slave_arready), //                                         .arready
		.hps_0_f2h_axi_slave_rid                        (mm_interconnect_0_hps_0_f2h_axi_slave_rid),     //                                         .rid
		.hps_0_f2h_axi_slave_rdata                      (mm_interconnect_0_hps_0_f2h_axi_slave_rdata),   //                                         .rdata
		.hps_0_f2h_axi_slave_rresp                      (mm_interconnect_0_hps_0_f2h_axi_slave_rresp),   //                                         .rresp
		.hps_0_f2h_axi_slave_rlast                      (mm_interconnect_0_hps_0_f2h_axi_slave_rlast),   //                                         .rlast
		.hps_0_f2h_axi_slave_rvalid                     (mm_interconnect_0_hps_0_f2h_axi_slave_rvalid),  //                                         .rvalid
		.hps_0_f2h_axi_slave_rready                     (mm_interconnect_0_hps_0_f2h_axi_slave_rready),  //                                         .rready
		.ccd_pixel_clock_bridge_out_clk_clk             (ccd_pixel_clock_bridge_clk),                    //           ccd_pixel_clock_bridge_out_clk.clk
		.accel_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                // accel_0_reset_sink_reset_bridge_in_reset.reset
		.accel_0_avalon_master_address                  (accel_0_avalon_master_address),                 //                    accel_0_avalon_master.address
		.accel_0_avalon_master_waitrequest              (accel_0_avalon_master_waitrequest),             //                                         .waitrequest
		.accel_0_avalon_master_read                     (accel_0_avalon_master_read),                    //                                         .read
		.accel_0_avalon_master_readdata                 (accel_0_avalon_master_readdata),                //                                         .readdata
		.accel_0_avalon_master_write                    (accel_0_avalon_master_write),                   //                                         .write
		.accel_0_avalon_master_writedata                (accel_0_avalon_master_writedata)                //                                         .writedata
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.ccd_pixel_clock_bridge_out_clk_clk                          (ccd_pixel_clock_bridge_clk),                          //                        ccd_pixel_clock_bridge_out_clk.clk
		.avalon_img_writer_rgbgray_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                      // avalon_img_writer_rgbgray_reset_reset_bridge_in_reset.reset
		.avalon_img_writer_rgbgray_avalon_master_address             (avalon_img_writer_rgbgray_avalon_master_address),     //               avalon_img_writer_rgbgray_avalon_master.address
		.avalon_img_writer_rgbgray_avalon_master_waitrequest         (avalon_img_writer_rgbgray_avalon_master_waitrequest), //                                                      .waitrequest
		.avalon_img_writer_rgbgray_avalon_master_burstcount          (avalon_img_writer_rgbgray_avalon_master_burstcount),  //                                                      .burstcount
		.avalon_img_writer_rgbgray_avalon_master_byteenable          (avalon_img_writer_rgbgray_avalon_master_byteenable),  //                                                      .byteenable
		.avalon_img_writer_rgbgray_avalon_master_write               (avalon_img_writer_rgbgray_avalon_master_write),       //                                                      .write
		.avalon_img_writer_rgbgray_avalon_master_writedata           (avalon_img_writer_rgbgray_avalon_master_writedata),   //                                                      .writedata
		.hps_0_f2h_sdram1_data_address                               (mm_interconnect_1_hps_0_f2h_sdram1_data_address),     //                                 hps_0_f2h_sdram1_data.address
		.hps_0_f2h_sdram1_data_write                                 (mm_interconnect_1_hps_0_f2h_sdram1_data_write),       //                                                      .write
		.hps_0_f2h_sdram1_data_writedata                             (mm_interconnect_1_hps_0_f2h_sdram1_data_writedata),   //                                                      .writedata
		.hps_0_f2h_sdram1_data_burstcount                            (mm_interconnect_1_hps_0_f2h_sdram1_data_burstcount),  //                                                      .burstcount
		.hps_0_f2h_sdram1_data_byteenable                            (mm_interconnect_1_hps_0_f2h_sdram1_data_byteenable),  //                                                      .byteenable
		.hps_0_f2h_sdram1_data_waitrequest                           (mm_interconnect_1_hps_0_f2h_sdram1_data_waitrequest)  //                                                      .waitrequest
	);

	soc_system_mm_interconnect_2 mm_interconnect_2 (
		.hps_0_h2f_axi_master_awid                                   (hps_0_h2f_axi_master_awid),                                          //                                  hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                 (hps_0_h2f_axi_master_awaddr),                                        //                                                      .awaddr
		.hps_0_h2f_axi_master_awlen                                  (hps_0_h2f_axi_master_awlen),                                         //                                                      .awlen
		.hps_0_h2f_axi_master_awsize                                 (hps_0_h2f_axi_master_awsize),                                        //                                                      .awsize
		.hps_0_h2f_axi_master_awburst                                (hps_0_h2f_axi_master_awburst),                                       //                                                      .awburst
		.hps_0_h2f_axi_master_awlock                                 (hps_0_h2f_axi_master_awlock),                                        //                                                      .awlock
		.hps_0_h2f_axi_master_awcache                                (hps_0_h2f_axi_master_awcache),                                       //                                                      .awcache
		.hps_0_h2f_axi_master_awprot                                 (hps_0_h2f_axi_master_awprot),                                        //                                                      .awprot
		.hps_0_h2f_axi_master_awvalid                                (hps_0_h2f_axi_master_awvalid),                                       //                                                      .awvalid
		.hps_0_h2f_axi_master_awready                                (hps_0_h2f_axi_master_awready),                                       //                                                      .awready
		.hps_0_h2f_axi_master_wid                                    (hps_0_h2f_axi_master_wid),                                           //                                                      .wid
		.hps_0_h2f_axi_master_wdata                                  (hps_0_h2f_axi_master_wdata),                                         //                                                      .wdata
		.hps_0_h2f_axi_master_wstrb                                  (hps_0_h2f_axi_master_wstrb),                                         //                                                      .wstrb
		.hps_0_h2f_axi_master_wlast                                  (hps_0_h2f_axi_master_wlast),                                         //                                                      .wlast
		.hps_0_h2f_axi_master_wvalid                                 (hps_0_h2f_axi_master_wvalid),                                        //                                                      .wvalid
		.hps_0_h2f_axi_master_wready                                 (hps_0_h2f_axi_master_wready),                                        //                                                      .wready
		.hps_0_h2f_axi_master_bid                                    (hps_0_h2f_axi_master_bid),                                           //                                                      .bid
		.hps_0_h2f_axi_master_bresp                                  (hps_0_h2f_axi_master_bresp),                                         //                                                      .bresp
		.hps_0_h2f_axi_master_bvalid                                 (hps_0_h2f_axi_master_bvalid),                                        //                                                      .bvalid
		.hps_0_h2f_axi_master_bready                                 (hps_0_h2f_axi_master_bready),                                        //                                                      .bready
		.hps_0_h2f_axi_master_arid                                   (hps_0_h2f_axi_master_arid),                                          //                                                      .arid
		.hps_0_h2f_axi_master_araddr                                 (hps_0_h2f_axi_master_araddr),                                        //                                                      .araddr
		.hps_0_h2f_axi_master_arlen                                  (hps_0_h2f_axi_master_arlen),                                         //                                                      .arlen
		.hps_0_h2f_axi_master_arsize                                 (hps_0_h2f_axi_master_arsize),                                        //                                                      .arsize
		.hps_0_h2f_axi_master_arburst                                (hps_0_h2f_axi_master_arburst),                                       //                                                      .arburst
		.hps_0_h2f_axi_master_arlock                                 (hps_0_h2f_axi_master_arlock),                                        //                                                      .arlock
		.hps_0_h2f_axi_master_arcache                                (hps_0_h2f_axi_master_arcache),                                       //                                                      .arcache
		.hps_0_h2f_axi_master_arprot                                 (hps_0_h2f_axi_master_arprot),                                        //                                                      .arprot
		.hps_0_h2f_axi_master_arvalid                                (hps_0_h2f_axi_master_arvalid),                                       //                                                      .arvalid
		.hps_0_h2f_axi_master_arready                                (hps_0_h2f_axi_master_arready),                                       //                                                      .arready
		.hps_0_h2f_axi_master_rid                                    (hps_0_h2f_axi_master_rid),                                           //                                                      .rid
		.hps_0_h2f_axi_master_rdata                                  (hps_0_h2f_axi_master_rdata),                                         //                                                      .rdata
		.hps_0_h2f_axi_master_rresp                                  (hps_0_h2f_axi_master_rresp),                                         //                                                      .rresp
		.hps_0_h2f_axi_master_rlast                                  (hps_0_h2f_axi_master_rlast),                                         //                                                      .rlast
		.hps_0_h2f_axi_master_rvalid                                 (hps_0_h2f_axi_master_rvalid),                                        //                                                      .rvalid
		.hps_0_h2f_axi_master_rready                                 (hps_0_h2f_axi_master_rready),                                        //                                                      .rready
		.ccd_pixel_clock_bridge_out_clk_clk                          (ccd_pixel_clock_bridge_clk),                                         //                        ccd_pixel_clock_bridge_out_clk.clk
		.avalon_img_writer_rgbgray_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                     // avalon_img_writer_rgbgray_reset_reset_bridge_in_reset.reset
		.accel_0_avalon_slave_address                                (mm_interconnect_2_accel_0_avalon_slave_address),                     //                                  accel_0_avalon_slave.address
		.accel_0_avalon_slave_write                                  (mm_interconnect_2_accel_0_avalon_slave_write),                       //                                                      .write
		.accel_0_avalon_slave_read                                   (mm_interconnect_2_accel_0_avalon_slave_read),                        //                                                      .read
		.accel_0_avalon_slave_readdata                               (mm_interconnect_2_accel_0_avalon_slave_readdata),                    //                                                      .readdata
		.accel_0_avalon_slave_writedata                              (mm_interconnect_2_accel_0_avalon_slave_writedata),                   //                                                      .writedata
		.accel_0_avalon_slave_waitrequest                            (mm_interconnect_2_accel_0_avalon_slave_waitrequest),                 //                                                      .waitrequest
		.avalon_camera_0_s1_address                                  (mm_interconnect_2_avalon_camera_0_s1_address),                       //                                    avalon_camera_0_s1.address
		.avalon_camera_0_s1_write                                    (mm_interconnect_2_avalon_camera_0_s1_write),                         //                                                      .write
		.avalon_camera_0_s1_read                                     (mm_interconnect_2_avalon_camera_0_s1_read),                          //                                                      .read
		.avalon_camera_0_s1_readdata                                 (mm_interconnect_2_avalon_camera_0_s1_readdata),                      //                                                      .readdata
		.avalon_camera_0_s1_writedata                                (mm_interconnect_2_avalon_camera_0_s1_writedata),                     //                                                      .writedata
		.avalon_img_writer_rgbgray_avalon_slave_address              (mm_interconnect_2_avalon_img_writer_rgbgray_avalon_slave_address),   //                avalon_img_writer_rgbgray_avalon_slave.address
		.avalon_img_writer_rgbgray_avalon_slave_write                (mm_interconnect_2_avalon_img_writer_rgbgray_avalon_slave_write),     //                                                      .write
		.avalon_img_writer_rgbgray_avalon_slave_read                 (mm_interconnect_2_avalon_img_writer_rgbgray_avalon_slave_read),      //                                                      .read
		.avalon_img_writer_rgbgray_avalon_slave_readdata             (mm_interconnect_2_avalon_img_writer_rgbgray_avalon_slave_readdata),  //                                                      .readdata
		.avalon_img_writer_rgbgray_avalon_slave_writedata            (mm_interconnect_2_avalon_img_writer_rgbgray_avalon_slave_writedata)  //                                                      .writedata
	);

	soc_system_irq_mapper irq_mapper (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq0_irq)  //    sender.irq
	);

	soc_system_irq_mapper irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_0_h2f_reset_reset),         // reset_in0.reset
		.clk            (ccd_pixel_clock_bridge_clk),     //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	assign h2f_reset_reset_n = ~rst_controller_reset_out_reset;

endmodule
